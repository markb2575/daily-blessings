2024-8-31|Mesra 25 1740|The Departure of St.Bessarion the Great, Pope Macarius III, 114th Patriarch|Psalm 1|What was your favorite verse and why?||
2024-9-1|Mesra 26 1740|The Martyrdom of St. Moses (Moises), St. Agabius, the Soldier |Psalm 3|What was your favorite verse and why?||
2024-9-2|Mesra 27 1740|The Martyrdom of Sts. Benjamin and Sister Eudoxia, St.Mary, the Armenian|Matthew 1|How many generations are between Abraham and Christ?|What does the word Emmanuel mean?|
2024-9-3|Mesra 28 1740|The Commemoration of the Patriarchs: Abraham, Isaac, and Jacob|Matthew 2|How did the wise men know that the child was king?|What prophecy did Jesus make to Egypt?|
2024-9-4|Mesra 29 1740|The Martyrdom of Sts. Athanasius, the Bishop and his servants|Matthew 3|What is the most important thing that was done by all who came to be baptized by John?|'But who comes _ is _ from me which I am not worthy to carry _'|Explain how the Father, the Son, and the Holy Spirit appeared during the baptism of the Lord Jesus by John
2024-9-5|Mesra 30 1740|The Departure of Malachi, the Prophet|Matthew 4|What did the Lord Jesus say when Satan asked him to turn the stones into bread?||
2024-9-6|Nasi 1 1740|The Departure of St. Eutychus |Matthew 5:1-26|What is the blessing for merciful people?|What must you do before receiving the Holy Communion?|
2024-9-7|Nasi 2 1740|The Departure of St. Titus, the Apostle |Matthew 5:27-48|Write your favorite verse from this week and what it means to you.||
2024-9-8|Nasi 3 1740|The Commemoration of Archangel Raphael, The Martyrdom of Sts.Andrianus, and his companions|Matthew 6:1-15|How should we perform charitable deeds?|'But if you _ men their _, your heavenly Father will also _ you. But if you do not forgive men their trespasses, _ will your Father forgive your trespasses.'|
2024-9-9|Nasi 4 1740|The Departure of St. Poimen, the Hermit|Matthew 6:16-34|What do we have to do when we are fasting?|'But seek first the _ and His righteousness, and all these things shall be _ to you.'|
2024-9-10|Nasi 5 1740|The Departure of St. Barsoum, the 'Naked'|Matthew 7:1-12|Why should we not judge others?|'_, and it will be given to you; _, and you will find; _, and it will be opened to you.'|
2024-9-11|Tout 1 1741|The Nayrouz Feast (Coptic New Year), The Departure of St. Bartholomew the Apostle |Matthew 7:13-29|Should we follow the narrow or wide path? Why?|Why would Jesus tell us to depart from Him?|
2024-9-12|Tout 2 1741|The Martyrdom of St. John the Baptist|Matthew 8:1-17|What miracles did Jesus perform?|Why did Jesus marvel at the Centurion?|
2024-9-13|Tout 3 1741||Matthew 8:18-34|What did Jesus say about the dead?|Why were the disciples scared? What did Jesus do?|
2024-9-14|Tout 4 1741|The Departure of St. Verena|Matthew 9:1-17|Write your favorite verse from this week and what it means to you.||
2024-9-15|Tout 5 1741|The Martyrdom of St. Sophia|Matthew 9:18-38|What did the bleeding woman believe?|How did the Pharisees think Jesus performed the miracle of casting out demons?|
2024-9-16|Tout 6 1741|The Martyrdom of Isaiah the Prophet, Son of Amoz|Matthew 10:1-23|Where did Jesus want to disciples to preach?|What did Jesus tell the disciples to do if they were turned away from a house or city?|
2024-9-17|Tout 7 1741|The Departure of Pope Dioscorus, 25th Pope of Alexandria|Matthew 10:24-42|'Therefore whoever _ Me before men, him I will also confess before My _ who is in _'|Who should we love first?|
2024-9-18|Tout 8 1741|The Departure of Moses the Prophet, The Martyrdom of Zacharias the Priest|Matthew 11:1-15|What did Jesus tell John's followers to tell him?||
2024-9-19|Tout 9 1741|The Martyrdom of St.Pisora the Bishop|Matthew 11:16-30|When should we thank our Father in heaven?|'Come to Me, all you who _ and are heavy _, and I will give you _'|
2024-9-20|Tout 10 1741|The Martyrdom of Sts. Youannes the Egyptian and his companions|Matthew 12:1-24|Does God want us to offer sacrifices? |What did Jesus say about the law of the Sabbath?|
2024-9-21|Tout 11 1741||Matthew 12:25-50|Write your favorite verse and what it means to you.||
2024-9-22|Tout 12 1741|The Commemoration of Archangel Michael|Matthew 13:1-15|Why did Jesus speak in parables?||
2024-9-23|Tout 13 1741||Matthew 13:16-33|What will happen to those who receive seeds on good ground?|How many parables did Jesus tell?|
2024-9-24|Tout 14 1741||Matthew 13:34-58|Jesus compares the kingdom of heaven to?|'So it will be at the end of the age. The _ will come forth, separate the _ from among the _, and cast them into the _ of fire.'|Where was Jesus rejected from?
2024-9-25|Tout 15 1741|The Translocation of the Body of St. Stephen the Archdeacon|Matthew 14:1-21|Who did King Herod think Jesus was?|How did Jesus feed the five thousand people?|
2024-9-26|Tout 16 1741||Matthew 14:22-36|Why do you think Jesus told the disciples to not be afraid?|Why did Peter begin to sink?|
2024-9-27|Tout 17 1741|The Feast of the Cross (Three days)|Matthew 15:1-20|What will happen if the blind lead the blind people?|Who did Jesus say are the blind people? Why?|
2024-9-28|Tout 18 1741|The Feast of the Cross (Three days)|Matthew 15:21-39|Write your favorite verse and what it means to you.||
2024-9-29|Tout 19 1741|The Feast of the Cross (Three days)|Matthew 16:1-12|When Jesus talked about bread to the disciples, what was He really talking about?||
2024-9-30|Tout 20 1741|The Departure of St. Theopista|Matthew 16:13-28|Who did Simon Peter say that Jesus is?|What did Jesus reveal to Peter after he said these things?|If anyone desires to come after Me, let him _ himself, and take up his _, and _ Me.'
2024-10-1|Tout 21 1741|The Commemoration of the Virgin St.Mary, the Theotokos, The Martyrdom of St. Cyprian the Bishop and St. Justina|Matthew 17:1-13|Who saw Jesus' transfiguration?|Jesus told the disciples not to speak of what they saw until?|
2024-10-2|Tout 22 1741||Matthew 17:14-27|Why were the disciples not able to cast out demons?|If you have _ as a _, you will say to this mountain, '_ from here to there'|
2024-10-3|Tout 23 1741||Matthew 18:1-20|Why does Jesus say we should become little children?|What will happen if we are lost like sheep?|
2024-10-4|Tout 24 1741|The Departure of St. Gregory, the Theologian|Matthew 18:21-35|When Jesus said to forgive your brother up to seventy times, what did He mean?|'So My heavenly Father also will do to you if each of you, from his _, does not_ his brother his _'|
2024-10-5|Tout 25 1741|The Departure of Jonah, the Great Prophet|Matthew 19:1-15|Write your favorite verse and what it means to you.||
2024-10-6|Tout 26 1741|The Annunciation of Zacharias the Priest with the Birth John the Baptist|Matthew 19:16-30|What did the rich man ask Jesus? How did He respond?|What does verse 30 mean?|
2024-10-7|Tout 27 1741||Matthew 20:1-16|What was the purpose of the story of the landowner and the laborers?|'So the last will be _, and the first _ For many are _, but few _'|
2024-10-8|Tout 28 1741||Matthew 20:17-34|What did Jesus tell his disciples?|What did the mother of Zebedee's son ask Jesus?|What does it mean to be last among others?
2024-10-9|Tout 29 1741||Matthew 21:1-22|What were people doing in the temple?|Why did Jesus condemns the fig tree?|
2024-10-10|Tout 30 1741||Matthew 21:23-46|Who believed the words of John the Baptist?|'The stone which the builder _ has become the chief _'|Who will receive the kingdom of heaven?
2024-10-11|Baba 1 1741|The Martyrdom of St. Anastasia|Matthew 22:1-22|From the parable: Why did the king throw out the man who was not dressed for the wedding?||
2024-10-12|Baba 2 1741||Matthew 22:23-46|Write your favorite verse and what it means to you.||
2024-10-13|Baba 3 1741|The Departure of Empress Theodora|Matthew 23:1-22|Did the Pharisees practice what they preached?||
2024-10-14|Baba 4 1741||Matthew 23:23-39|What is Jesus warning the Pharisee about?|What does it mean that the Pharisee drink from a cup clean on the outside, but dirty on the inside? |
2024-10-15|Baba 5 1741|The Martyrdom of St. Paul, Patriarch of Constantinople|Matthew 24:1-14|What will happen to those who follow Christ at the end?|Why should we continue to trust in the Lord?|
2024-10-16|Baba 6 1741|The Departure of the Righteous Hannah, Mother of Samuel, the Prophet|Matthew 24:15-31|'And He will send His _ with a great sound of a _, and they will gather together His elect from the four _, from one end of heaven to the other'||
2024-10-17|Baba 7 1741|The Departure of St. Paul of Tammoh|Matthew 24:32-51|Why must we always be ready?||
2024-10-18|Baba 8 1741||Matthew 25:1-23|What happened to the five foolish women?|What did the servants with five and two talents do with them?|
2024-10-19|Baba 9 1741||Matthew 25:24-46|Write your favorite verse and what it means to you.||
2024-10-20|Baba 10 1741||Matthew 26:1-25|What did Jesus say the woman anointing His feet was doing?|How did the disciples know Judas was going to betray Jesus?|
2024-10-21|Baba 11 1741|The Departure of St. James, Patriarch of Antioch |Matthew 26:26-46|What did this Passover meal with Jesus represent?|Where did Jesus go to pray at night?|What were the disciples doing while Jesus was praying?
2024-10-22|Baba 12 1741|The Commemoration of the Honorable Archangel Michael, The Martyrdom of St. Matthew the Evangelist|Matthew 26:47-68|When the disciple cut the ear of the servant, what did Jesus say?|Who was the high priest who Jesus saw at night?|
2024-10-23|Baba 13 1741|The Departure of St. Zacharias, the Monk|Matthew 26:69-75|What did Peter do outside the courtyard?|What did he do after?|
2024-10-24|Baba 14 1741|The Departure of St. Philip, One of the Seven Deacons |Matthew 27:1-14|What is the Field of Blood?|What did Jesus say in front of Pilate?|
2024-10-25|Baba 15 1741|The Martyrdom of St. Panteleimon, the Physician|Matthew 27:15-31|Who did Pilate release instead of Jesus?|What did the Roman soldiers do with Jesus?|
2024-10-26|Baba 16 1741||Matthew 27:32-48|Write your favorite verse and what it means to you.||
2024-10-27|Baba 17 1741|The Departure of St. Dioscorus II, 31st Pope of Alexandria |Matthew 27:49-66|After Jesus yielded His spirit, what happened?|Whose tomb was Jesus buried in?|What were the Pharisees afraid the disciples would do?
2024-10-28|Baba 18 1741||Matthew 28|What did the angel tell the women who were walking to Jesus' tomb?|What did the chief priests pay the soldiers to say?|Go therefore and make _ of all the nations, _ them in the name of the _ and of the _ and of the _'
2024-10-29|Baba 19 1741||Exodus 1|What happened to the Hebrews after a new Pharoh came to rule?|What did this new King do with the Hebrew babies that were born?|
2024-10-30|Baba 20 1741|The Departure of the Great St. John Colobos (the Short) |Exodus 2|What did the Levite woman who had a son do with him?|What happened to Moses when he fled Egypt?|
2024-10-31|Baba 21 1741|The Commemoration of the Theotokos, the Virgin St. Mary, The Departure of Joel the Prophet|Exodus 3|What was the name of the mountain on which the Lord appeared to Moses from the burning bush?|When Moses asked what he should say when the Egyptians ask 'What is his name?'?|
2024-11-1|Baba 22 1741|The Martyrdom of St. Luke the Evangelist|Exodus 4:1-13|What happened when Moses threw the staff on the ground?|Why did Moses not want to go to Egypt?|
2024-11-2|Baba 23 1741||Exodus 4:14-31|Write your favorite verse and what it means to you.||
2024-11-3|Baba 24 1741||Exodus 5|What did Pharoh do when Moses and Aaron asked to let His people go?|Who did the Isrealites blame when their work became harder?|
2024-11-4|Baba 25 1741||Exodus 6:1-13|'I will free you from being _ to them, and I will redeem you with an outstretched arm and with _ acts of _  I will take you as my own people, and I will be your God. Then you will know that I am the Lord your God, who brought you out from under the yoke of the _'||
2024-11-5|Baba 26 1741|The Martyrdom of St. Timon the Apostle|Psalm 8|What was your favorite verse and why?||
2024-11-6|Baba 27 1741|The Martyrdom of St. Macarius, Bishop of Edko |Exodus 7:1-13|What was the first miracle Moses and Aaron performed?|What did Pharoh do in response?|
2024-11-7|Baba 28 1741|Martyrdom of the Sts. Marcian and Mercurius |Exodus 7:14-25|What was the first plague performed?|What happened to the Egyptians because of this?|
2024-11-8|Baba 29 1741|The Martyrdom of St. Demetrius of Thessalonica|Exodus 8:1-19|What was the second plague? The third?|Why did Pharoh not listen?|
2024-11-9|Baba 30 1741||Exodus 8:20-32|Write your favorite verse and what it means to you.||
2024-11-10|Hatour 1 1741|The Martyrdom of St. Cleopas the Apostle, one of the two Disciples of Emmaus|Exodus 9:1-12|What was the fifth and sixth plague?||
2024-11-11|Hatour 2 1741||Exodus 9:13-35|What was the seventh plague?|What did Pharoh do after this plague? Did he let this Isrealites go?|
2024-11-12|Hatour 3 1741|The Martyrdom of St. Athanasius and His sister, Irene, St. Aghathon|Exodus 10:1-11|What did God say the next plague was going to be?||
2024-11-13|Hatour 4 1741|The Martyrdom of Sts. John and James, Bishops of Persia|Exodus 10:12-29|What was the ninth plague?|What did Pharoh allow the Isrealites to do?|
2024-11-14|Hatour 5 1741|The Martyrdom of St. Timothy, the Deacon|Exodus 11|Why was their going to be a great cry in Egypt?||
2024-11-15|Hatour 6 1741||Exodus 12:1-20|What did the Isrealites need to do to be saved from the strike of the firstborns?||
2024-11-16|Hatour 7 1741|The Martyrdom of St. George, the Alexandrian |Exodus 12:21-36|Write your favorite verse and what it means to you.||
2024-11-17|Hatour 8 1741||Exodus 12:37-51|Why did the Isrealites take the bread unleavened?|What happened to the Isrealites this Passover?|
2024-11-18|Hatour 9 1741|The Assembly of the First Ecumenical Council at Nicea|Exodus 13|How many days will the eat unleavened bread?|What was leading this Isrealites through the wilderness?|
2024-11-19|Hatour 10 1741|The Martyrdom of the Fifty Virgins and their mother St. Sophia|Exodus 14:1-14|Who was behind the Isrealites when they reached the Red Sea?|What did Moses tell those who were scared?|
2024-11-20|Hatour 11 1741|The Departure of St. Anna (Hannah), the mother of the Holy Virgin St. Mary |Exodus 14:15-31|What stood between the Isrealites and the Egyptians?|What happened after the Isrealites crossed on dry land?|
2024-11-21|Hatour 12 1741||Exodus 15:1-13|'I will sing to the Lord, For He has _ gloriously! The horse and its _ He has thrown into the _!'||
2024-11-22|Hatour 13 1741||Exodus 15:14-27|Why was the water undrinkable for the Isrealites?|What did Moses do to satisfy their thirst?|
2024-11-23|Hatour 14 1741||Exodus 16:1-21|Write your favorite verse and what it means to you.||
2024-11-24|Hatour 15 1741|The Martyrdom of St. Mari-Mina, the Wonder Worker|Exodus 16:22-36|What happened to the bread that the people kept for the morning after?||
2024-11-25|Hatour 16 1741|Start of The Holy Nativity Fast|Exodus 17|What did Moses do when the people said they were thirsty?|How did the Isrealites win against the Amaleks?|
2024-11-26|Hatour 17 1741|The Departure of St. John Chrysostom |Exodus 18:1-12|What did Jethro do when he rejoiced for the Isrealites being released from Egypt?||
2024-11-27|Hatour 18 1741|The Martyrdom of St. Philip the Apostle |Exodus 18:13-27|When Moses was judging the people, why did Jethro say this was wrong?|What did Moses do to help this issue?|
2024-11-28|Hatour 19 1741||Exodus 19|How long have the Isrealites been in the wilderness at this point?|Why was it that only Moses and Aaron could travel up Mount Sinai?|
2024-11-29|Hatour 20 1741||Exodus 20|What is the first comandment given to Moses? The fifth?|'Do not fear; for God has come to _ you, and that His _may be before you, so that you may not _'|
2024-11-30|Hatour 21 1741|The Commemoration of the Virgin St. Mary, the Theotokos, The Departure of St. Gregory, the Wonder Worker|Exodus 21:1-17|Write your favorite verse and what it means to you.||
2024-12-1|Hatour 22 1741||Exodus 21:18-36|List some verses that state a sin and the punishment? |Do you think the death punishments are a literal death, or have another meaning?|
2024-12-2|Hatour 23 1741|The Departure of St. Cornelius the Centurion|Exodus 22:1-14|What is the punishment for those who steal? |What does it mean to make restitution?|
2024-12-3|Hatour 24 1741|The Commemoration of the Twenty-Four Presbyters|Exodus 22:15-30|What verse specifically mentions to not worship other gods? What are we told to not do when loaning people money (hint: verse 25)?|What are we told to not do when loaning people money (hint: verse 25)?|
2024-12-4|Hatour 25 1741|The Martyrdom of St. Mercurius Known as the Saint with the Two Swords|Exodus 23:1-19|What verse(s) is an example of the saying 'love your enemies?' ||
2024-12-5|Hatour 26 1741||Exodus 23:20-33|'You shall not bow down to their gods, nor _ them, nor do according to their _ ; but you shall utterly overthrow them and completely break down their sacred _'||
2024-12-6|Hatour 27 1741|The Martyrdom of St. James the Persian |Exodus 24|Who did God call to worship Him?|How long was Moses on the mountain?|
2024-12-7|Hatour 28 1741||Exodus 25:1-22|Write your favorite verse and what it means to you.||
2024-12-8|Hatour 29 1741|The Martyrdom of St. Catherine of Alexandria |Psalm 10|What was your favorite verse and why?||
2024-12-9|Hatour 30 1741|The Martyrdom of St. Macarius, Monk St. John El-Qalyuby|Exodus 26:1-14|What is surrounding the tabernacle?|What color(s) did God say it should be?|
2024-12-10|Kiahk 1 1741||Exodus 26:15-37|What wood is the tabernacle made of?|What is overlaid on the wood?|
2024-12-11|Kiahk 2 1741||Exodus 27|What meterial is used for the south side of the tabernacle?|Who watched over the lampstand so that it continuously burns?|
2024-12-12|Kiahk 3 1741|The Martyrdom of St. Bestavros, the New Martyr|Exodus 28:1-21|Who was chosen to be the priests?|What color(s) of thread should be used for the ephod?|
2024-12-13|Kiahk 4 1741|The Martyrdom of St. Andrew, One of the Twelve Apostles |Exodus 28:22-43|'So Aaron shall bear the names of the sons of Israel on the _ of judgment over his _, when he goes into the holy place, as a memorial before the Lord _'|What was engraved on the plate of gold?|
2024-12-14|Kiahk 5 1741||Exodus 29:1-21|Write your favorite verse and what it means to you.||
2024-12-15|Kiahk 6 1741||Exodus 29:22-46|What should be done with the ram after it has been consecrated?|What and when should be offered on the altar daily?|
2024-12-16|Kiahk 7 1741|The Departure of St. Mettaos El-Fakhoury (Matthew the Poor)|Exodus 30:1-16|What incense should be offered on the altar?|What should the Isrealites do as they are taking a census?|
2024-12-17|Kiahk 8 1741|The Martyrdom of St. Esi and His Sister Thecla, Two Saints: Barbara and Juliana|Exodus 30:17-38|What spices are used in annointing oil?||
2024-12-18|Kiahk 9 1741||Exodus 31|Why is the Sabbath, the seventh day, a day of rest?||
2024-12-19|Kiahk 10 1741||Exodus 32:1-14|When Moses was on the mountain a long time, what did the people ask Aaron to do?|When God was angry with the Isrealites, what did Moses do?|
2024-12-20|Kiahk 11 1741||Exodus 32:15-35|What did Moses do when he saw the people dancing?|What did Moses pray for? How did God respond?|
2024-12-21|Kiahk 12 1741|The Departure of St. John the Confessor|Exodus 33|Write your favorite verse and what it means to you.||
2024-12-22|Kiahk 13 1741|The Commemoration of the Honorable Archangel Raphael|Exodus 34:1-17|What did the Lord command Moses to do?||
2024-12-23|Kiahk 14 1741||Exodus 34:18-35|Why is the Feast of Unleavened Bread during the month of Abib?|What happened to Moses when he came down Mount Sinai?|
2024-12-24|Kiahk 15 1741|The Departure of St. Gregory Patriarch of the Armenians|Exodus 35:1-19|List some of the articles within the tabernacle?||
2024-12-25|Kiahk 16 1741|The Departure of the Righteous Gideon, One of the Judges of Israel|Exodus 35:20-35|What were some of the offerings people brought to the tabernacle?||
2024-12-26|Kiahk 17 1741||Psalm 25|What was your favorite verse and why?||
2024-12-27|Kiahk 18 1741||Psalm 26|What was your favorite verse and why?||
2024-12-28|Kiahk 19 1741||Exodus 37|Write your favorite verse and what it means to you.||
2024-12-29|Kiahk 20 1741|The Departure of Haggai the Prophet|Exodus 38:1-20|What was hanging on the West side of the tabernacle?||
2024-12-30|Kiahk 21 1741|The Commemoration of the Pure Virgin St.Mary, the Theotokos, The Martyrdom of St. Barnabas, One of the Seventy Apostles|Psalm 33|What was your favorite verse and why?||
2024-12-31|Kiahk 22 1741|The Commemoration of the Honorable Archangel Gabriel, the Announcer|Psalm 36|What was your favorite verse and why?||
2025-1-1|Kiahk 23 1741|The Departure of David, the Prophet and King, St. Timothy, the Anchorite|Exodus 40:1-21|What should Aaron and his son's do before entering the tabernacle?||
2025-1-2|Kiahk 24 1741|The Departure of St. Ignatius, Theophorus, Patriarch of Antioch|Exodus 40:22-38|Where was the lampstand placed?|When could the priest enter the tabernacle?|
2025-1-3|Kiahk 25 1741||Psalm 40|What was your favorite verse and why?||
2025-1-4|Kiahk 26 1741|The Martyrdom of St. Anastasia|James 1|Write your favorite verse and what it means to you.||
2025-1-5|Kiahk 27 1741||James 2|What does James mean when he says we should not have faith with partiality?|'For judgment is without _ to the one who has shown _ Mercy _ over judgment'|
2025-1-6|Kiahk 28 1741|The Holy Nativity Fast|James 3|What does this verse mean, 'But no man can tame the tongue. It is an unruly evil, full of deadly poison. With it we bless our God and Father, and with it we curse men, who have been made in the similtude of God.'|What is James saying we should be careful of becoming? Why?|
2025-1-7|Kiahk 29 1741|The Holy Nativity Feast|James 4|What does God resist? What does He give to the humble?|James tells us that tomorrow is not guaranteed. What does he compare our lives to?|
2025-1-8|Kiahk 30 1741||James 5|'You also be _ Establish your _, for the coming of the Lord is at _'|What should we do if someone is suffering? Cheeful? Sick?|
2025-1-9|Toba 1 1741|The Martyrdom of St. Stephen the Archdeacon|Psalm 84|What was your favorite verse and why?||
2025-1-10|Toba 2 1741||Psalm 95|What was your favorite verse and why?||
2025-1-11|Toba 3 1741|The Martyrdom of the Children of Bethlehem |Psalm 96|What was your favorite verse and why?||
2025-1-12|Toba 4 1741|The Departure of St. John the Evangelist |Psalm 98|What was your favorite verse and why?||
2025-1-13|Toba 5 1741||Joshua 1|What did the Lord tell Joshua he will do for him? (hint: the Lord said he did the same thing with Moses)|Did the people obey the Lord's commands, which were told by Joshua?|
2025-1-14|Toba 6 1741|The Circumcision Feast|Joshua 2|How did Rahab help the two men from Acacia Grove?|What did Rahab request from the men in return for helping them?|
2025-1-15|Toba 7 1741||Joshua 3|Where did Joshua and the children of Israel travel to?|What happened to the 12 men that were chosen from each tribe?|
2025-1-16|Toba 8 1741||Joshua 4|What is the significance of the stones that were moved to the lodging place?|What happened to the Jordan waters once the priests stepped on land?|
2025-1-17|Toba 9 1741||Joshua 5|What did the Lord command to Joshua in regards to circumcision?|What did the commander of the army of the Lord tell Joshua at the end of the chapter?|
2025-1-18|Toba 10 1741|Paramouni of the Honorable Theophany Feast (Epiphany)|Joshua 6:1-25|Write your favorite verse and what it means to you.||
2025-1-19|Toba 11 1741|The Holy Epiphany (Baptism of the Lord Christ)|Joshua 7|What happened to Achan as his punishment?||
2025-1-20|Toba 12 1741|The Second day of the feast of Holy Theophany, Commemoration of the Honorable Archangel Michael|Joshua 8:1-25|'And it will be, when you have _ the city, that you shall set the city on _'|What happened to the king of Ai|
2025-1-21|Toba 13 1741|Feast of the Wedding of Cana of Galilee, Martyrdom of St.Demiana|Joshua 9|What did the inhabitants of Gibeon do when they heard about Joshua and what happened at Jericho and Ai?|What was their punishment for lying about their identity?|
2025-1-22|Toba 14 1741||Joshua 10:1-27|What natural disaster took place that killed the Amorites?|What happened to the five kings?|
2025-1-23|Toba 15 1741|The Departure of Obadiah, the Prophet|Joshua 11|Why did the city of Hazor get burned?|Who were the only people that made peace with the children of Israel?|
2025-1-24|Toba 16 1741|The Martyrdom of St.Philotheus|Joshua 12|How many kings total did Joshua and the children of Israel conquer on the west side of the Jordan?||
2025-1-25|Toba 17 1741||Joshua 13: 1-23|Write your favorite verse and what it means to you.||
2025-1-26|Toba 18 1741|The Departure of St.James, Bishop of Nisibis|Joshua 14|What was the only thing the Levites recieved?|What did Caleb do during the time of Moses?|
2025-1-27|Toba 19 1741||Joshua 15: 1-19|What did Caleb state was the condition to recieve his daughter, Achsah?|Who took Caleb's daughter?|
2025-1-28|Toba 20 1741||Joshua 16|Where did the Canaanites dwell?||
2025-1-29|Toba 21 1741|The Departure of the Virgin St.Mary, the Mother of God, St.Hilaria the daughter of Emperor Zeno|Joshua 17|What did the children of Israel do to the Canaanites in an attempt to drive them out?|What did Joshua tell the children of Joseph in response to them stating they have little land?|
2025-1-30|Toba 22 1741|The Departure of the Great St.Anba Anthony the Father of all Monks|Joshua 18|How many tribes did not recieve their inheritance when the children of Israel gathered at Shiloh?|What did Joshua command from the men in terms of recieving land?|
2025-1-31|Toba 23 1741|The Martyrdom of St.Timothy the Apostle|Joshua 19:1-22|'The inheritance of the children of _ was included in the share of the children of _, for the share of the children of _ was too much for them.'|What land did the children of Issachar recieve?|
2025-2-1|Toba 24 1741|The Departure of St.Mary the Ascetic|Joshua 20|What was your favorite verse and why?||
2025-2-2|Toba 25 1741||Joshua 21:1-26|'And the children of _ gave these cities with their common-lands by lot to the _, as the _ had commanded by the hand of _'||
2025-2-3|Toba 26 1741||Joshua 22:1-29|What did Joshua say about where to return as the Lord had promised?|'Far be it from us that we should _ against the Lord, and turn from _ the Lord this day, to build an _ for burnt offerings, for _ offerings or for _ , besides the altar of the Lord our God which is before his _'|
2025-2-4|Toba 27 1741|The Commemoration of the Honorable Archangel Suriel|Joshua 23|What did Joshua tell the people in his farewell address?|What does Joshua state will happen if the people turn from God to serve others?|
2025-2-5|Toba 28 1741||Joshua 24:1-29|But Joshua said to the people 'You cannot _ the Lord, for he is a _ God. He is a _ God; he will not forgive your _ nor your _''|How old was Joshua when he died?|
2025-2-6|Toba 29 1741|The Departure of St.Eksanie |Psalm 103|What was your favorite verse and why?||
2025-2-7|Toba 30 1741||Psalm 111|What was your favorite verse and why?||
2025-2-8|Amshir 1 1741|The Commemoration of the Second Universal Council in the city of Constantinople|Acts 1:1-11|Write your favorite verse and what it means to you.||
2025-2-9|Amshir 2 1741|The Departure of the Great St.Anba Paul, the First Hermit|Acts 1:12-26|What did the eleven disciples do before making a decision about another person for their ministry?|Who was chosen to replace Judas as disciple?|
2025-2-10|Amshir 3 1741|Jonah's (Nineveh) Fast, The Departure of St.James the Monk|Acts 2:1-21|What happened on the day of Pentecost?|Filled with the Holy Spirit, what were the disciples able to do?|
2025-2-11|Amshir 4 1741|Jonah's (Nineveh) Fast|Acts 2:22-47|After preaching, what did Peter do with those listening?|About how many people were baptized that day?|
2025-2-12|Amshir 5 1741|Jonah's (Nineveh) Fast|Acts 3|Instead of alms, what did St.Peter do for the lame man?|When people were amazed by this miracle, what did Peter say to them?|
2025-2-13|Amshir 6 1741|Jonah's (Nineveh) Feast|Acts 4:1-17|What happened to Peter and John after this miracle?|When the Sanhedrin asked Peter by what power has he performed this miracle, how did he respond?|
2025-2-14|Amshir 7 1741||Acts 4:18-37|Once Peter and John were released they prayed to the Lord, 'grant to Your _ that with all boldness they may _ Your word, by stretching out Your _ to heal, and that signs and _ may be done through the name of Your holy Servant _'||
2025-2-15|Amshir 8 1741|Presentation of the Lord into the Temple, Departure of St.Simeon the Elder|Acts 5:1-16|Write your favorite verse and what it means to you.||
2025-2-16|Amshir 9 1741||Acts 5:17-42|What happened when the apostles were locked in prison? Where did they go after?|Why were the captain and officers afraid of arresting the apostles?|
2025-2-17|Amshir 10 1741||Acts 6|What did the false witnesses claim St. Stephen taught about Jesus and the Temple?|'And it shall come to pass that whoever _ on the name of the _ shall be _'|
2025-2-18|Amshir 11 1741||Acts 7:1-22|What was the covenant God gave to Abraham?|Which Holy Forefather begot the twelve patriarchs ?|
2025-2-19|Amshir 12 1741|The Commemoration of the Honorable Archangel Michael |Acts 7:23-43|How many years did Moses stay in the land of Midian?|What did the Jewish people do in the wilderness after they were released from Egypt?|
2025-2-20|Amshir 13 1741||Acts 7:44-60|How was St.Stephen martyred?|'Look! I see the _ opened and the Son of Man _ at the right hand of _!'|
2025-2-21|Amshir 14 1741|The Departure of St.Severus, Patriarch of Antioch|Acts 8:1-25|What happened while Philip was preaching in Samaria?|What did Peter say to Simon when he tried to buy power with money?|
2025-2-22|Amshir 15 1741||Acts 8:26-40|Write your favorite verse and what it means to you.||
2025-2-23|Amshir 16 1741|The Departure of St.Elizabeth, Mother of St.John the Baptist|Acts 9:1-25|Who spoke to Saul on his journey to Damascus? What did He say?|'Go, for he is a _ of Mine to bear My name before _, kings, and the children of _’'|
2025-2-24|Amshir 17 1741|Start of Holy Great Fast, The Martyrdom of St.Mina the Monk|Acts 9:26-43|Who brought Saul to the Apostles?|What happened to Tabitha? What did Peter do?|
2025-2-25|Amshir 18 1741||Acts 10:1-23|What was Cornelius' job?|During Peter's vison he heard a voice? What did it say the first and second time?|
2025-2-26|Amshir 19 1741||Acts 10:24-46|What did Cornelius do when St. Peter entered his house?|While Peter was preaching to the household and friends of Cornelius, something unusual happened. What was it that happened?|
2025-2-27|Amshir 20 1741||Acts 11:1-15|'Then the _ told me to go with them,_ Moreover these six brethren accompanied me, and we entered the man’s house.'|The Church in Jerusalem sent which individual to Antioch?|
2025-2-28|Amshir 21 1741|The Commemoration of the Virgin St.Mary, the Theotokos|Acts 11:16-30|'When they heard these things they became silent; and they _ God, saying, ‘Then God has also _ to the Gentiles _ to life.’'|Where were the disciples first called Christians?|
2025-3-1|Amshir 22 1741||Acts 12|Write your favorite verse and what it means to you.||
2025-3-2|Amshir 23 1741||Acts 13:1-12|Where did Paul and Barnabas travel to?|Who was traveling with Barnabas and Saul ?|
2025-3-3|Amshir 24 1741|The Martyrdom of St.Timothy and St.Matthias|Acts 13:13-35|What happened at Antioch of Pesidia ?|How many nations did God destroy in Canaan for his people ?|
2025-3-4|Amshir 25 1741|The Martyrdom of Sts.Philemon, Apphia, and their son Archippus|Acts 13:36-52|You will not allow Your Holy One to see corruption' a prophecy was said about?|What did the people seek after hearing to St. Paul ?|
2025-3-5|Amshir 26 1741|The Departure of the Righteous Hosea, the Prophet|Acts 14:1-13|Who believed in Iconium ?|What did the people at Lystra do when they saw the miracle ?|
2025-3-6|Amshir 27 1741|The Departure of St.Eustathius, Patriarch of Antioch|Acts 14:14-28|Where did the apostles go after the stoning ?|What did they do on ther way back to Lystra, Antioch and Iconium ?|
2025-3-7|Amshir 28 1741||Acts 15:1-21|What did the people of Judea teach the others brethren ?|'So God, who knows the _, acknowledged them by giving them the _, just as He did to us, and made no distinction between us and them, _ their hearts by_'|
2025-3-8|Amshir 29 1741||Acts 15:22-41|Write your favorite verse and what it means to you.||
2025-3-9|Amshir 30 1741||Acts 16:1-20|What did St. Paul do to St. Timothy before they left ?|What led St. Paul to believe that the Lord was calling him to preach in Macedonia?|
2025-3-10|Baramhat 1 1741|The Martyrdom of St.Alexandrus, the Soldier|Acts 16:21-40|How did St. Paul and St. Silas exceedingly trouble the city?|How many members of the Philippian jailer’s household were baptized?|
2025-3-11|Baramhat 2 1741||Acts 17:1-15|St. Paul explained and proved that two things were necessary for the Christ to do. What were they?||
2025-3-12|Baramhat 3 1741||Acts 17:16-34|Where did the philosophers take St. Paul to hear him speak about his 'new doctrine?'|Paul found one particular altar in Athens, What was the inscription on this altar?|
2025-3-13|Baramhat 4 1741||Acts 18:1-11|Why were Aquila and Priscilla in Corinth?|Which ruler of the synagogue in Corinth became a Christian with his household?|
2025-3-14|Baramhat 5 1741||Acts 18:12-28|Which ruler of the synagogue in Corinth became a Christian with his household?|Which ruler of the synagogue in Corinth became a Christian with his household?|
2025-3-15|Baramhat 6 1741|The Martyrdom of St.Dioscorus|Acts 19:1-22|Write your favorite verse and what it means to you.||
2025-3-16|Baramhat 7 1741|The Martyrdom of St.Mary the Israelite|Acts 19:23-41|What did the silversmiths cry out?|What crime did the city clerk of Ephesus convict Gaius and Aristarchus?|
2025-3-17|Baramhat 8 1741|The Martyrdom of St.Matthias, the apostle|Psalm 134|What was your favorite verse and why?||
2025-3-18|Baramhat 9 1741||Psalm 136|What was your favorite verse and why?||
2025-3-19|Baramhat 10 1741|The Feast of the Cross|Psalm 141|What was your favorite verse and why?||
2025-3-20|Baramhat 11 1741|The Martyrdom of St.Basil the Bishop|Esther 1|What caused King Ahasuerus to become angry?|What did the King do in response?|
2025-3-21|Baramhat 12 1741|Commemoration of the Honorable Archangel Michael|Esther 2|What is Esther's other name? Why did she hide her people?|What did Bigthan and Teresh try to do? What happened to them instead?|
2025-3-22|Baramhat 13 1741|The Martyrdom of the Forty Martyrs of Sebaste|Esther 3|Write your favorite verse and what it means to you.||
2025-3-23|Baramhat 14 1741||Esther 4|What would happen if a person went before the king without being called?|What did Esther ask of the Jewish people?|
2025-3-24|Baramhat 15 1741|The Departure of St.Sarah the Nun|Esther 5|What request did Esther make of the king?|What was Haman's plan for Mordecai?|
2025-3-25|Baramhat 16 1741||Esther 6|When the king could not sleep he read some records. What did he find?|To honor Mordecai, what did King Ahasuerus do?|
2025-3-26|Baramhat 17 1741|The Departure of Lazarus, the beloved of the Lord, The Martyrdom of St.Sidhom Bishay in Domiat|Esther 7|What did Queen Esther say at the second banquet?|What happened to Haman in the end?|
2025-3-27|Baramhat 18 1741||Esther 8|Why did Queen Esther cry in front of the king?|What was the new decree that was signed by the king?|
2025-3-28|Baramhat 19 1741||Esther 9:1-17|What happened to the Jews on the thirteenth day of themonth of Adar?|What occured on the fourteenth day of the month of Adar?|
2025-3-29|Baramhat 20 1741||Esther 9:18-32|Write your favorite verse and what it means to you.||
2025-3-30|Baramhat 21 1741|The Commemoration of the Theotokos, the Pure Virgin St.Mary, The Martyrdom of Sts.Theodore and Timothy|Esther 10|What position did Mordecai have with the king?||
2025-3-31|Baramhat 22 1741||Psalm 143|What was your favorite verse and why?||
2025-4-1|Baramhat 23 1741|The Departure of the Great Prophet Daniel|Psalm 144|What was your favorite verse and why?||
2025-4-2|Baramhat 24 1741||Ruth 1|After Naomi's sons had passed away, what did her daughter-in-laws do? What about Ruth?|Where did Naomi and Ruth travel to?|
2025-4-3|Baramhat 25 1741||Ruth 2|What did Naomi ask Ruth to do?|Blessed be he of the _ , who has not forsaken His _ to the _ and the _!' Why does Naomi rejoice?|
2025-4-4|Baramhat 26 1741|The Departure of St.Euphrasia, the Virgin|Ruth 4:13-22|Who are the descendants of Ruth and Boaz?||
2025-4-5|Baramhat 27 1741|The Commemoration of the Crucifixion of our Lord Jesus Christ, The Departure of St.Macarius the Great|Psalm146|What was your favorite verse and why?||
2025-4-6|Baramhat 28 1741|The Departure of Emperor Constantine the Great|Psalm 147|What was your favorite verse and why?||
2025-4-7|Baramhat 29 1741|Annunciation Feast, The Commemoration of the Resurrection of the Lord Christ from the dead|Psalm 148|What was your favorite verse and why?||
2025-4-8|Baramhat 30 1741|The Commemoration of Archangel Gabriel the Announcer, The Departure of Samson, One of the Judges of Israel|Psalm 150|What was your favorite verse and why?||
2025-4-9|Baramouda 1 1741|The Departure of St.Silvanus the monk, Aaron the priest|1 Samuel 1:1-18|What was the vow that Hannah made to the Lord?|What did Eli the priest think of Hannah?|
2025-4-10|Baramouda 2 1741|The Martyrdom of St.Christopher|1 Samuel 1:19-28|What did Hannah bring up with her to offer to the Lord?|'For this child I _, and the Lord _ me my petition which I asked of Him'|
2025-4-11|Baramouda 3 1741||1 Samuel 2:1-17|'No one is holy like the _, For there is none besides You, Nor is there any _ like our God.'|After Elkanah went to his house,who did Samuel stay with?|
2025-4-12|Baramouda 4 1741|Lazarus Saturday|1 Samuel 2:18-36|Write your favorite verse and what it means to you.||
2025-4-13|Baramouda 5 1741|Entry of our Lord into Jerusalem (Hosanna Sunday)||||
2025-4-14|Baramunda 6 1741|Holy Pascha||||
2025-4-15|Baramouda 7 1741|Holy Pascha||||
2025-4-16|Baramunda 8 1741|Holy Pascha||||
2025-4-17|Baramouda 9 1741|Covenant Thursday||||
2025-4-18|Baramouda 10 1741|Good Friday||||
2025-4-19|Baramouda 11 1741|||||
2025-4-20|Baramouda 12 1741|Glorious Feast of the Resurrection||||
2025-4-21|Baramouda 13 1741||1 Samuel 3|What did Eli tell Samuel to say when the Lord calls him?|Why was God upset with Eli?|
2025-4-22|Baramouda 14 1741||1 Samuel 4|What happened to the ark of God during battle?|What happened to Eli when he heard that the ark of God was captured?|
2025-4-23|Baramouda 15 1741||1 Samuel 5|What happened to Dagon when the ark of God was placed in the house of Dagon?|What did the Philistines decide to do with the ark of God?|
2025-4-24|Baramouda 16 1741|The Martyrdom of St.Antipas, Bishop of Pergamos|1 Samuel 6|What did the priests tell the Philistines to do when they are sending the ark of God to its place?|How did the people of Shemesh celebrate the return of the ark of God?|
2025-4-25|Baramouda 17 1741|The Martyrdom of St.James One of the Twelve Apostles, Brother of St.John the Beloved, The Departure of St.Nicodemus|1 Samuel 7|What did the children of Israel do after Samuel spoke to them?|What did God do when the Philistines came near to battle the children of Israel?|
2025-4-26|Baramouda 18 1741||1 Samuel 8|Write your favorite verse and what it means to you.||
2025-4-27|Baramouda 19 1741|Thomas’ Sunday|1 Samuel 9:1-14|What did Kish ask of his son Saul?|What did Saul ask the young women who were going out to draw water?|
2025-4-28|Baramouda 20 1741||1 Samuel 9:15-27|Who said 'I am the Seer'?|'But as for your donkeys that were lost three days ago, do not be _ about them, for they have been _'|
2025-4-29|Baramouda 21 1741|The Commemoration of the Virgin St.Mary, the Theotokos|1 Samuel 10:1-16|'Then the _ of the Lord will come upon you and you will _ with them and be turned into another _'||
2025-4-30|Baramouda 22 1741||1 Samuel 10:17-27|'I brought up Israel out of _, and delivered you from the hand of the _ and from the hand of all _ and from those who oppressed you.'|Who was appointed a king over the people of Israel?|
2025-5-1|Baramouda 23 1741|The Martyrdom of St.George Prince of the Martyrs|1 Samuel 11|How many children of Israel and how many men of Judah went out with Saul?|What did the people do to Saul in Gilgal?|
2025-5-2|Baramouda 24 1741||1 Samuel 12|Why did the people of Israel cry out to the Lord?|'So Samuel called to the Lord, and the Lord sent _ and _that day.'|
2025-5-3|Baramouda 25 1741||1 Samuel 13|Write your favorite verse and what it means to you.||
2025-5-4|Baramouda 26 1741|The Martyrdom of St.Sonos|1 Samuel 14:1-25|What is the name of Saul’s son?|'But if they say thus ‘Come up to us, then we will go up. For the Lord has _ them into our hand, and this will be a sign to us.'|
2025-5-5|Baramouda 27 1741||1 Samuel 14:26-52|Why were the people not able to eat from the honey?||
2025-5-6|Baramouda 28 1741|The Martyrdom of St.Milius, the Ascetic|1 Samuel 15:1-16|God told Saul to go attack who?|Why was God upset with Saul?|
2025-5-7|Baramouda 29 1741|The Departure of St.Erastus, the Apostle|1 Samuel 15:17-35|What was Saul planning to do with the sheep and oxen ?|How does Saul feel about not obeying God’s commandment?|
2025-5-8|Baramouda 30 1741|Martyrdom of St. Mark the Evangelist|1 Samuel 16|'You shall _for Me the one I _ to you.'|Why did Saul send messengers to Jesse?|
2025-5-9|Bashans 1 1741|The Nativity of the Blessed Virgin Mary the Mother of God|1 Samuel 17:1-20|Who said 'why have you come out to line up for battle?'|How many brothers did David have?|
2025-5-10|Bashans 2 1741|The Departure of the Righteous Job|1 Samuel 17:21-39|Write your favorite verse and what it means to you.||
2025-5-11|Bashans 3 1741|The Departure of St.Jason, One of the Seventy Disciples|1 Samuel 17:40-58|Why did David take off the sword and the armor?|What two things did David use to defeat Goliath?|
2025-5-12|Bashans 4 1741||1 Samuel 18:1-16|What did Jonathan give to David?|Who said 'Saul has slain his thousands, and David his ten thousands'.|
2025-5-13|Bashans 5 1741|The Martyrdom of Jeremiah the Prophet|1 Samuel 18:17-30|What is the name of Saul’s daughter that David married?|'And Saul was still more _of David. So Saul became _’s enemy continually.'|
2025-5-14|Bashans 6 1741||1 Samuel 19|Who warned David that Saul wants to kill him?|What did Michal tell Saul’s messengers when they went to take David?|
2025-5-15|Bashans 7 1741||1 Samuel 20:1-21|Who said the following to David? 'By no means! You shall not die!'|Where did David hide?|
2025-5-16|Bashans 8 1741|The Commemoration of the Ascension of Our Lord jesus Christ in Heaven, The Martyrdom of St.John of Senhout|1 Samuel 20:22-42|'But the lad did not know anything. Only _ and _ knew of the matter.'|Why did David and Jonathan cry?|
2025-5-17|Bashans 9 1741|The Departure of St.Helena, the Queen|1 Samuel 21|Write your favorite verse and what it means to you.||
2025-5-18|Bashans 10 1741|The Departure of the Three Holy Young Men Hananiah, Azariah, and Mishael|1 Samuel 22|How many men were with David?|Who told David that Saul had killed the Lord's priests?|
2025-5-19|Bashans 11 1741||1 Samuel 23:1-13|Who said the following verse? 'God has delivered him into my hand, for he has shut himself in by entering a town that has gates and bars.'|Where did David escape from?|
2025-5-20|Bashans 12 1741|The Commemoration of the Honorable Archangel Michael|1 Samuel 23:14-29|David and his men were in the Wilderness of Maon, in the plain on the south of|What did they call the place after Saul returned from pursuing David?|
2025-5-21|Bashans 13 1741|The Departure of St.Arsenius, the Tutor of the Emperor's Children|1 Samuel 24|What did David do to Saul while Saul was in the cave?|'May the Lord _ you with _ for what you have done to me this day.'|
2025-5-22|Bashans 14 1741||1 Samuel 25:1-20|What was the name of the very rich man?|Who was going to give David and his men bread, wine, sheep, grain, and cakes of figs?|
2025-5-23|Bashans 15 1741|The Martyrdom of St.Simon the Zealot (Simon the Canaanite), one of the Twelve Apostles, 400 martyrs in Dandara|1 Samuel 25:21-44|Who was holding a feast in his house?|'But Saul had given _ his daughter, David’s _, to Palti the son of Laish, who was from _'|
2025-5-24|Bashans 16 1741||1 Samuel 26|Write your favorite verse and what it means to you.||
2025-5-25|Bashans 17 1741|The Departure of St.Epiphanius, Bishop of Cyprus|1 Samuel 27|Who was David trying to escape from?|How long did David dwell in the country of the Philistines?|
2025-5-26|Bashans 18 1741|The Commemoration of the feast of Pentecost|1 Samuel 28|Who did the Philistines want to have a war against?|Who said the following: 'Therefore I have called you, that you may reveal to me what I should do.'|
2025-5-27|Bashans 19 1741||1 Samuel 29|Then the Princes of the _said, 'what are these _doing here?'|'As soon as you are up early in the _and have _, depart.'|
2025-5-28|Bashans 20 1741||1 Samuel 30:1-15|What did David and his men find when they returned to Ziklag?|What did David and his men do to the Egyptian that they found in the field?|
2025-5-29|Bashans 21 1741|The Holy Feast of Ascension|1 Samuel 30:16-31|'Now when David came to Ziklag, he sent some of the _ to the elders of _'|'Those who were in _, and to all the places where David himself and his _ were accustomed to rove.'|
2025-5-30|Bashans 22 1741|The Departure of St.Andronicus, one of the Seventy Disciples|1 Samuel 31|Who killed Saul’s three sons?|What did the inhabitants of Jabesh Gilead do when they heard what the Philistines had done to Saul?|
2025-5-31|Bashans 23 1741|The Departure of St.Junia, One of the Seventy Disciples|2 Samuel 1:1-12|Write your favorite verse and what it means to you.||
2025-6-1|Bashans 24 1741|Entry of the Lord into Egypt|2 Samuel 1:13-27|What did David do to the man who killed Saul?|They were swifter than _they were stronger than _' **|
2025-6-2|Bashans 25 1741||2 Samuel 2:1-16|Where did God tell David to go?|What was the name of Saul’s son who reigned as king over Israel?|
2025-6-3|Bashans 26 1741|The Martyrdom of St.Thomas the Apostle|2 Samuel 2:17-32|Whose servants won the battle?|Then Abner called to Joab and said, shall the _devour forever'? **|
2025-6-4|Bashans 27 1741|The Departure of Lazarus the Beloved of the Lord|2 Samuel 3:1-20|How many sons were born to David in Hebron?|For the Lord has spoken of David, saying ‘By the hand of David I will _ My people Israel from the hand of the _ and the hand of all their _' **|
2025-6-5|Bashans 28 1741||2 Samuel 3:21-39|Who did Joab kill?|How did King David feel when he found out that Abner is dead?|
2025-6-6|Bashans 29 1741|The Departure of St.Simon the Stylite|2 Samuel 4|What is the name of Jonathan’s son who was lame in his feet?|What did David command his men to do with the head of Ishbosheth?|
2025-6-7|Bashans 30 1741||2 Samuel 5|Write your favorite verse and what it means to you.||
2025-6-8|Paona 1 1741|The Holy Pentecost Feast|2 Samuel 6|Why did God strike Uzzah?|Why did king David decide to go bring the ark of God from the house of Obed-Edom to the City of David?|
2025-6-9|Paona 2 1741|Start of The Apostles' Fast|2 Samuel 7:1-17|What is the name of the prophet that King David spoke to and said 'See now, I dwell in a house of cedar, but the ark of God dwells inside tent curtains'?||
2025-6-10|Paona 3 1741||2 Samuel 7:18-29|Now, O Lord God, the word which You have spoken concerning Your _ and concerning his _, establish it forever and do as You have said.' **|And now, O Lord God, You are God, and Your words are _, and You have promised this goodness to Your _' **|
2025-6-11|Paona 4 1741||2 Samuel 8|What did David take from  Hadadezer the son of Rehob?|So David reigned over all Israel; and David administered _ and _ to all his people.' **|
2025-6-12|Paona 5 1741|The Departure of St.James the Oriental, the Confessor, The Martyrdom of St.Bifam|2 Samuel 9|What was the name of the servant from the house of Saul?|Do not fear, for I will surely show you _ for _ your father’s sake, and will restore to you all the _ of Saul your grandfather.' **|
2025-6-13|Paona 6 1741|The Martyrdom of St.Theodore, the Monk|2 Samuel 10|What did Hanun do to David’s servants?|And when all the kings who were servants to _saw that they were defeated by Israel, they made _ with Israel and served them.' **|
2025-6-14|Paona 7 1741||2 Samuel 11:1-11|Write your favorite verse and what it means to you.||
2025-6-15|Paona 8 1741||2 Samuel 11:12-27|Why did king David want Joab to put Uriah in the forefront of the hottest battle?|What happened to Uriah the Hittitie during the war?|
2025-6-16|Paona 9 1741|The Departure of Samuel the Prophet|2 Samuel 12:1-15|Who was the prophet that God sent to David?|What did the prohet say would happen because of David's sin?|
2025-6-17|Paona 10 1741||2 Samuel 12:16-31|What did King David do when he found out?|Then he took their king’s _ from his head. Its weight was a talent of gold, with precious stones. And it was set on _ head.' **|
2025-6-18|Paona 11 1741|The Martyrdom of St.Claudius|2 Samuel 13:1-20|What is the name of Absalom’s sister?|So that the hatred with which he hated her was greater than the _ with which he had loved her' **|
2025-6-19|Paona 12 1741|The Commemoration of Archangel Michael, The Departure of St.Euphemia|2 Samuel 13:21-39|What did Absalom do to Amnon?|How long was Absalom at Geshur?|
2025-6-20|Paona 13 1741|The Commemoration of the Archangel Gabriel, the Announcer|2 Samuel 14:1-14|And when the woman of _ spoke to the king, she fell on her face to the ground and _ herself, and said, 'Help, O _ !' **|What did the woman of Tekoa pretend that her problem was?|
2025-6-21|Paona 14 1741||2 Samuel 14:15-33|Write your favorite verse and what it means to you.||
2025-6-22|Paona 15 1741||2 Samuel 15:1-16|As soon as you hear the sound of the _, then you shall say, _ reigns in Hebron!’ ' **|Who did king David flee from?|
2025-6-23|Paona 16 1741|The Departure of Abba Nofer the Anchorite|2 Samuel 15:17-37|How many men followed king David from Gath?|What did king David ask Hushai the Archite to do?|
2025-6-24|Paona 17 1741|The Departure of St.Latsoun el-Bahnasawy|2 Samuel 16|What did Ziba bring to king David?|Did Ahithophel give good or bad advice?|
2025-6-25|Paona 18 1741||2 Samuel 17:1-14|Who did Ahithophel and Absalom want to kill?|Did Hushai agree with Ahithophel’s advice?|
2025-6-26|Paona 19 1741||2 Samuel 17:15-29|Arise and cross over the _ quickly. For thus has Ahithophel advised _ you.' **|What did Ahithophel do when he saw that his advice was not followed?|
2025-6-27|Paona 20 1741|The Departure of Elisha, the Prophet|2 Samuel 18:1-18|What did king David command Joab, Abishai, and Ittai regarding Absalom?|What did they do with Absalom after he died?|
2025-6-28|Paona 21 1741||2 Samuel 18:19-32|Write your favorite verse and what it means to you.||
2025-6-29|Paona 22 1741||2 Samuel 19:1-20|Now therefore, arise, go out and speak _ to your servants. For I swear by the Lord, if you do not go out, not one will stay with you this _' **|Did king David want to kill Shimei?|
2025-6-30|Paona 23 1741|The Departure of St.Abba Nouub the Confessor|2 Samuel 19:21-43|Did Brazillai agree to go across the Jordan with king David?|We have ten _ in the king; therefore we also have more _ to David than you.' **|
2025-7-1|Paona 24 1741|The Martyrdom of the Mighty Saint Abba Moses the Ethiopian|2 Samuel 20|And the king took the ten women, his _ whom he had left to keep the house, and put them in _ and supported them' **|What were the names of the two priests of Israel?|
2025-7-2|Paona 25 1741||2 Samuel 21|How long was the famine and why did it occur?|How many giants did the Philistines have? What happened to them?|
2025-7-3|Paona 26 1741||2 Samuel 22:1-25|The Lord is my _ and my fortress and my deliverer; The God of my _, in whom I will trust; My shield and the horn of my _' **||
2025-7-4|Paona 27 1741|The Martyrdom of St.Ananias, the Apostle|2 Samuel 22:26-51|What does verse 29-31 mean to you?|What is King David doing in the last 5 verses?|
2025-7-5|Paona 28 1741||2 Samuel 23:1-19|Write your favorite verse and what it means to you.||
2025-7-6|Paona 29 1741|The Martyrdom of the Seven Ascetics in Tounah Mount|Psalm 17|What was your favorite verse and why?||
2025-7-7|Paona 30 1741|The Nativity of St.John, the Baptist|2 Samuel 24:1-13|What did God ask King David to do?|What were the three options that the prophet Gad gave to David from God?|
2025-7-8|Abib 1 1741|The Martyrdom of St.Febronia, the Ascetic|2 Samuel 24:14-25|Which of the three happened to Israel?|What did David do to withdraw the plague on Israel?|
2025-7-9|Abib 2 1741|The Departure of St.Jude, the Apostle|Daniel 1|How many sons did Judah have and what were their names?|What happened after the 10 days when Daniel told the steward to test his servants?|
2025-7-10|Abib 3 1741||Daniel 2:1-23|What caused the king to be angry and commanded that all the wise men of Babylon be killed?|How was the kings secret revealed to Daniel?|
2025-7-11|Abib 4 1741||Daniel 2:24-49|Describe Daniel's vision of the secret.|How did king Nebuchadnezzar react to Daniel’s vision?|
2025-7-12|Abib 5 1741|The Apostles' Feast (Martyrdom of St. Peter & St. Paul)|Daniel 3:1-15|Write your favorite verse and what it means to you.||
2025-7-13|Abib 6 1741|The Martyrdom of St.Theodosia and her companions|Daniel 3:16-30|Who was the fourth man that the king saw in the firery furnace with Shadrach, Meshach, and Abed-Nego?||
2025-7-14|Abib 7 1741|The Departure of St.Shenouda, the Archimandrite|Daniel 4:1-18|Explain the vision that king Nebuchadnezzar saw in his dream.|What did he ask Daniel (Belteshazzar) to do?|
2025-7-15|Abib 8 1741||Daniel 4:19-37|What advice did Daniel give the king after telling him the interpretation of his dream?|At the end of the chapter, did king Nebuchadnezzar praise God?|
2025-7-16|Abib 9 1741|The Martyrdom of St.Simon son of Clopas, the Apostle and Bishop of Jerusalem|Daniel 5:1-12|What was the reward that the king Belshazzar would grant to whoever interpreted the writing?|The queen, because of the words of the king and his lords, came to the banquet hall. The queen spoke, saying, ‘_! Do not let your thoughts _ you, nor let your _change.' **|
2025-7-17|Abib 10 1741|The Martyrdom of St.Theordore, Bishop of Pentapolis|Daniel 5:13-31|Why did the king want Daniel to interpret the writing?|What was the interpretation for the word TEKEL?|
2025-7-18|Abib 11 1741|The Martyrdom of Sts.John and Simon, his cousin|Daniel 6:1-17|All the governors of the kingdom, the administrators and satraps, the counselors and advisors, have consulted together to establish a _ and to make a firm _, that whoever _any god or man for thirty days, except you, O king, shall be cast into the _' **|Why did king Damaris put Daniel into the lions’ den?|
2025-7-19|Abib 12 1741|The Commemoration of Archangel Michael|Daniel 6:18-28|Write your favorite verse and what it means to you.||
2025-7-20|Abib 13 1741||Daniel 7:1-14|How many beasts did Daniel see in his vision?|Describe each of the beasts.|
2025-7-21|Abib 14 1741|The Martyrdom of St.Proconius of Jerusalem|Daniel 7:15-28|What was the first interpretation of the four beasts in Daniel’s vision?|What was the true interpretation of the four beasts in Daniel’s vision?|
2025-7-22|Abib 15 1741|The Departure of St.Ephrem the Syrian|Daniel 8:1-14|Describe the two animals that Daniel saw in his vision.||
2025-7-23|Abib 16 1741|The Departure of St.John, the Owner of the Golden Gospel|Daniel 8:15-27|What did Gabriel say this vision represents?|What nations did the animals represent?|
2025-7-24|Abib 17 1741|The Martyrdom of St.Euphemia|Daniel 9|What did you learn from the humility of Daniel's prayer?||
2025-7-25|Abib 18 1741|The Martyrdom of St.James the Apostle, the Brother of the Lord, Bishop of Jerusalem|Psalm 63|What was your favorite verse and why?||
2025-7-26|Abib 19 1741||Psalm 64|Write your favorite verse and what it means to you.||
2025-7-27|Abib 20 1741|The Martyrdom of St.Theordore of Shotep|Daniel 10|Which angel is mentioned in Daniel's vision? They are reffered to as 'one of the chief princes'.||
2025-7-28|Abib 21 1741|The Commemoration of the Lady, the Virgin St.Mary|Psalm 75|What was your favorite verse and why?||
2025-7-29|Abib 22 1741||Psalm 76|What was your favorite verse and why?||
2025-7-30|Abib 23 1741|The Martyrdom of St.Longinus the Soldier, St.Marina of Antioch|Mark 1:1-20|Who is the messenger who God sent in front of Jesus Christ to prepare His path?|On the Epiphany day the Holy Trinity appeared. How did the Father appear? The son? The Holy Spirit?|
2025-7-31|Abib 24 1741||Mark 1:21-45|Why did Lord Jesus Christ not let the demons speak?|What happened when our Lord Jesus Christ breathed His last?|
2025-8-1|Abib 25 1741|The Martyrdom of St.Isaac, St.Hilaria|Mark 2:1-12|What did the friends of the paralytic man do to reach Jesus Christ ?|Why were the people angry from what our Lord said ?|
2025-8-2|Abib 26 1741|The Departure of the Upright St.Joseph, the Carpenter|Mark 2:13-28|Write your favorite verse and what it means to you.||
2025-8-3|Abib 27 1741|The Martyrdom of St.Apamon |Mark 3:1-19|What were the Pharisee's reaction to this miracle?|'For He _ many, so that as many as had afflictions pressed into Him about _'|
2025-8-4|Abib 28 1741|The Departure of St.Mary Magdalene|Mark 3:20-35|'If a kingdom is divided against itself, _'|What is the only sin that will have no forgiveness?|
2025-8-5|Abib 29 1741||Mark 4:1-20|What happened to the seed that fell on the wayside? The stony ground? Among thorns? On good ground?|'_ they may see and not perceive, and _ They may and not understand. Lest they should turn and their _'|
2025-8-6|Abib 30 1741|The Martyrdom of Sts.Mercurius and Ephraem|Mark 4:21-41|Our Lord Jesus Christ said that the Kingdom of God is like?|What did our Lord Jesus say to the disciples ?|
2025-8-7|Mesra 1 1741|Start of St. Mary's Fast|Mark 5:1-20|What happened to the herd of swine when the unclean spirits entered them ?|What did our Lord Jesus say to the demon, possessed man when he begged Him to leave him?|
2025-8-8|Mesra 2 1741|The Departure of St.Paesa (Athanasia)|Mark 5:21-43|The sick woman had a strong faith, because she said?|Which disciples were taken to Jairus' house?|
2025-8-9|Mesra 3 1741||Mark 6:1-13|Write your favorite verse and what it means to you.||
2025-8-10|Mesra 4 1741|The Departure of Hezekiah, the Righteous King|Mark 6:14-29|Why did King Heord arrest St.John the Baptist?|What did Herodia's daughter ask Herod for? Did he accept or refuse?|
2025-8-11|Mesra 5 1741|The Martyrdom of St.John the Soldier|Mark 6:30-44|'And Jesus when He came out, saw a _ and was moved with compassion for them because they were like _ Not having a _'|How many baskets were left over?|
2025-8-12|Mesra 6 1741|The Martyrdom of St.Julietta, The Departure of St.Jacob al-Baradai|Mark 6:45-56|How did Jesus appear to the disciples?|What was the blind man's name?|
2025-8-13|Mesra 7 1741||Mark 7:1-23|'These people honor me with their _, but their _ is far from me.'|Write a verse about honoring your father and mother.|
2025-8-14|Mesra 8 1741||Mark 7:24-37|Who was the woman who approached Jesus? What did she ask of Him?|Our Lord Jesus Christ made the deaf _ and _ speak.|
2025-8-15|Mesra 9 1741||Mark 8:1-21|What did the Pharisees asked our Lord Jesus Christ?|When Jesus warned His disciples of the Pharisee's and Herod, what did they think He was talking about?|
2025-8-16|Mesra 10 1741|The Martyrdom of St.Pihebs, St.Matra|Mark 8:22-38|Write your favorite verse and what it means to you.||
2025-8-17|Mesra 11 1741|The Departure of St.Moisis, Bishop of Ouseem|Mark 9:1-13|Who did Jesus take on the mountain with Him? What happened?|Who will come before the second coming?|
2025-8-18|Mesra 12 1741|The Commemoration of the Honorable Archangel Michael|Mark 9:14-32|What did Our Lord Jesus Christ see when He came down form the mountain?|'If you can believe , _ are possible to him who believes.'|
2025-8-19|Mesra 13 1741|Transfiguration Feast|Mark 9:33-50|'For whoever gives you a _ to drink in _ because you belong to Christ, assuredly, I say to you, he will by no means lose his _'|'Have salt in yourselves and have _'|
2025-8-20|Mesra 14 1741||Mark 10:1-16|Why can a man not divorce his wife?|What did Jesus say about children?|
2025-8-21|Mesra 15 1741||Mark 10:17-31|Based on what Jesus said, how do we get to heaven? List three points.|'Children, how hard it is for those who _ to enter the kingdom of God!'|
2025-8-22|Mesra 16 1741|Assumption of St. Mary's Body|Mark 10:32-52|'But whoever desires to become great among you shall be your _ and whoever of you desires to be _ shall be slave of all. For even the Son of Man did not come to be served, but to _ and to give His _ a ransom for many.'||
2025-8-23|Mesra 17 1741|The Martyrdom of St.James the Soldier|Mark 11:1-14|Write your favorite verse and what it means to you.||
2025-8-24|Mesra 18 1741|The Departure of St.Alexander, Patriarch of Constantinople|Mark 11:15-33|Why was Jesus angry? Write the verse below.|'And whenever you stand praying, if you have anything _ anyone, _ him, that your Father in heaven may also forgive you your _'|
2025-8-25|Mesra 19 1741||Mark 12:1-17|The stone which the builders rejected, has become the _|'Render to _ the things that are Caesar’s, and to God the things that are _'|
2025-8-26|Mesra 20 1741|The Martyrdom of the Seven Young Men of Ephesus|Mark 12:18-34|'When we rise from the death we will be like _ in heaven.'|'He is not the God of the _, but the God of the _'|
2025-8-27|Mesra 21 1741|The Commemoration of the Virgin St.Mary, the Mother of God, The Departure of St.Irene|Mark 12:35-44|‘The Lord said to my _, 'Sit at My right hand, Till I make Your _ Your footstool.''|Who said this prophesy?|
2025-8-28|Mesra 22 1741|The Departure of Micah, the Prophet, St.Augustine|Mark 13:1-22|What the prophecy that our Lord Jesus Christ said about the temple ?|'But when they arrest you and deliver you up, _ beforehand, or premeditate what you will speak. But whatever is given you in that hour, speak that; for it is not you who _, but the _'|
2025-8-29|Mesra 23 1741||Mark 13:23-37|'Heaven and earth will pass away, but My _ will by no means _'|Who is the only one who knows the hour and day?|
2025-8-30|Mesra 24 1741||Mark 14:1-16|Write your favorite verse and what it means to you.||
2025-8-31|Mesra 25 1741|The Departure of St.Bessarion, the Great|Mark 14:17-31|What did Jesus tell His disciples during Passover Feast?|What did Jesus say will happen after the ressurection?|
2025-9-1|Mesra 26 1741|The Martyrdom of St.Moses and his Sister Sarah|Mark 14:32-52|Where did they go after the last supper?|What sign did Judas give to arrest Jesus?|
2025-9-2|Mesra 27 1741|The Martyrdom of Sts.Benjamin and his Sister Eudoxia, St.Mary the Armenian|Mark 14:53-72|When Jesus said 'I am' what did the high priest do?|What did St.Peter do when he realized he had denied Jesus?|
2025-9-3|Mesra 28 1741|The Commemoration of the Patriarchs: Abraham, Issac, and Jacob|Mark 15:1-20|What did Pilate ask our Lord Jesus Christ?|What was Pilate's tradition on the feast? Who did he release?|
2025-9-4|Mesra 29 1741|The Martyrdom of Sts. Athanasius, the Bishop and his servants|Mark 15:21-47|What is the name of the man who helped carry the cross with Jesus?|What happened when Jesus Christ breathed His last?|
2025-9-5|Mesra 30 1741|The Departure of Malachi, the Prophet|Mark 16|Who went to the tomb early in the morning?|'Go into all the world and preach the _ to every creature. He who believes and is _ will be _ ; but he who does not believe will be _'|